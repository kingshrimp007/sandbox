module vc_outbufs # (
    parameter D_WIDTH = 32,
    parameter VID_BITS = 6,
    parameter PORTS = 5,
    parameter CHANNELS = 12,
    localparam NUM_REQ = PORTS * CHANNELS
) (
    
);


endmodule