module sym_butterfly_wrapper #(
    parameter integer PORTS = 64
) (
    input logic clk,
    input logic 
);
